package Def ;

typedef 5 L;
typedef 4 EXTEST ;
typedef 2 SAMPLE_PRELOAD ;
typedef 31 BYPASS ;
typedef 17 DBA  ;
typedef 16 DTM ;
typedef 1 IDCODE ;

endpackage